LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity zeroCheck_tb is
end zeroCheck_tb;

architecture behavioral of zeroCheck is

component zeroCheck

port(
    input:      in std_logic_vector(7 downto 0);
    output:     out std_logic--_vector(7 downto 0)
);
end component;

signal inpt: std_logic_vector(7 downto 0);
signal otpt: std_logic;--_vector(7 downto 0);

begin

z1: zeroCheck port map(input=>inpt,output=>otpt);

process

type pattern_type is record

inpt: std_logic_vector (7 downto 0);

otpt: std_logic;--_vector (7 downto 0);

end record;

type pattern_array is array (natural range <>) of pattern_type;

constant patterns : pattern_array :=
(
("00000000",'1'),
("00000001",'0'),
("00000010",'0'),
("00000011",'0'),
("00000100",'0'),
("00000101",'0'),
("00000110",'0'),
("00000111",'0'),
("00001000",'0'),
("00001001",'0'),
("00001010",'0'),
("00001011",'0'),
("00001100",'0'),
("00001101",'0'),
("00001110",'0'),
("00001111",'0'),
("00010000",'0'),
("00010001",'0'),
("00010010",'0'),
("00010011",'0'),
("00010100",'0'),
("00010101",'0'),
("00010110",'0'),
("00010111",'0'),
("00011000",'0'),
("00011001",'0'),
("00011010",'0'),
("00011011",'0'),
("00011100",'0'),
("00011101",'0'),
("00011110",'0'),
("00011111",'0'),
("00100000",'0'),
("00100001",'0'),
("00100010",'0'),
("00100011",'0'),
("00100100",'0'),
("00100101",'0'),
("00100110",'0'),
("00100111",'0'),
("00101000",'0'),
("00101001",'0'),
("00101010",'0'),
("00101011",'0'),
("00101100",'0'),
("00101101",'0'),
("00101110",'0'),
("00101111",'0'),
("00110000",'0'),
("00110001",'0'),
("00110010",'0'),
("00110011",'0'),
("00110100",'0'),
("00110101",'0'),
("00110110",'0'),
("00110111",'0'),
("00111000",'0'),
("00111001",'0'),
("00111010",'0'),
("00111011",'0'),
("00111100",'0'),
("00111101",'0'),
("00111110",'0'),
("00111111",'0'),
("01000000",'0'),
("01000001",'0'),
("01000010",'0'),
("01000011",'0'),
("01000100",'0'),
("01000101",'0'),
("01000110",'0'),
("01000111",'0'),
("01001000",'0'),
("01001001",'0'),
("01001010",'0'),
("01001011",'0'),
("01001100",'0'),
("01001101",'0'),
("01001110",'0'),
("01001111",'0'),
("01010000",'0'),
("01010001",'0'),
("01010010",'0'),
("01010011",'0'),
("01010100",'0'),
("01010101",'0'),
("01010110",'0'),
("01010111",'0'),
("01011000",'0'),
("01011001",'0'),
("01011010",'0'),
("01011011",'0'),
("01011100",'0'),
("01011101",'0'),
("01011110",'0'),
("01011111",'0'),
("01100000",'0'),
("01100001",'0'),
("01100010",'0'),
("01100011",'0'),
("01100100",'0'),
("01100101",'0'),
("01100110",'0'),
("01100111",'0'),
("01101000",'0'),
("01101001",'0'),
("01101010",'0'),
("01101011",'0'),
("01101100",'0'),
("01101101",'0'),
("01101110",'0'),
("01101111",'0'),
("01110000",'0'),
("01110001",'0'),
("01110010",'0'),
("01110011",'0'),
("01110100",'0'),
("01110101",'0'),
("01110110",'0'),
("01110111",'0'),
("01111000",'0'),
("01111001",'0'),
("01111010",'0'),
("01111011",'0'),
("01111100",'0'),
("01111101",'0'),
("01111110",'0'),
("01111111",'0'),
("10000000",'0'),
("10000001",'0'),
("10000010",'0'),
("10000011",'0'),
("10000100",'0'),
("10000101",'0'),
("10000110",'0'),
("10000111",'0'),
("10001000",'0'),
("10001001",'0'),
("10001010",'0'),
("10001011",'0'),
("10001100",'0'),
("10001101",'0'),
("10001110",'0'),
("10001111",'0'),
("10010000",'0'),
("10010001",'0'),
("10010010",'0'),
("10010011",'0'),
("10010100",'0'),
("10010101",'0'),
("10010110",'0'),
("10010111",'0'),
("10011000",'0'),
("10011001",'0'),
("10011010",'0'),
("10011011",'0'),
("10011100",'0'),
("10011101",'0'),
("10011110",'0'),
("10011111",'0'),
("10100000",'0'),
("10100001",'0'),
("10100010",'0'),
("10100011",'0'),
("10100100",'0'),
("10100101",'0'),
("10100110",'0'),
("10100111",'0'),
("10101000",'0'),
("10101001",'0'),
("10101010",'0'),
("10101011",'0'),
("10101100",'0'),
("10101101",'0'),
("10101110",'0'),
("10101111",'0'),
("10110000",'0'),
("10110001",'0'),
("10110010",'0'),
("10110011",'0'),
("10110100",'0'),
("10110101",'0'),
("10110110",'0'),
("10110111",'0'),
("10111000",'0'),
("10111001",'0'),
("10111010",'0'),
("10111011",'0'),
("10111100",'0'),
("10111101",'0'),
("10111110",'0'),
("10111111",'0'),
("11000000",'0'),
("11000001",'0'),
("11000010",'0'),
("11000011",'0'),
("11000100",'0'),
("11000101",'0'),
("11000110",'0'),
("11000111",'0'),
("11001000",'0'),
("11001001",'0'),
("11001010",'0'),
("11001011",'0'),
("11001100",'0'),
("11001101",'0'),
("11001110",'0'),
("11001111",'0'),
("11010000",'0'),
("11010001",'0'),
("11010010",'0'),
("11010011",'0'),
("11010100",'0'),
("11010101",'0'),
("11010110",'0'),
("11010111",'0'),
("11011000",'0'),
("11011001",'0'),
("11011010",'0'),
("11011011",'0'),
("11011100",'0'),
("11011101",'0'),
("11011110",'0'),
("11011111",'0'),
("11100000",'0'),
("11100001",'0'),
("11100010",'0'),
("11100011",'0'),
("11100100",'0'),
("11100101",'0'),
("11100110",'0'),
("11100111",'0'),
("11101000",'0'),
("11101001",'0'),
("11101010",'0'),
("11101011",'0'),
("11101100",'0'),
("11101101",'0'),
("11101110",'0'),
("11101111",'0'),
("11110000",'0'),
("11110001",'0'),
("11110010",'0'),
("11110011",'0'),
("11110100",'0'),
("11110101",'0'),
("11110110",'0'),
("11110111",'0'),
("11111000",'0'),
("11111001",'0'),
("11111010",'0'),
("11111011",'0'),
("11111100",'0'),
("11111101",'0'),
("11111110",'0')

);
begin

for n in patterns'range loop

inpt <= patterns(n).inpt;

wait for 1 ns;

assert otpt = patterns(n).otpt
report "bad output value" severity error;
end loop;
assert false report "end of test" severity note;

wait;
end process;
end behavioral;